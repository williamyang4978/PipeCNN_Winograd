// mult_add_fix8bx16bx4.v

// Generated using ACDS version 18.0.1 261

`timescale 1 ps / 1 ps
module mult_add_fix8bx16bx4 (
		input  wire        clock0,  //  clock0.clock0
		input  wire [15:0] dataa_0, // dataa_0.dataa_0
		input  wire [15:0] dataa_1, // dataa_1.dataa_1
		input  wire [15:0] dataa_2, // dataa_2.dataa_2
		input  wire [15:0] dataa_3, // dataa_3.dataa_3
		input  wire [7:0]  datab_0, // datab_0.datab_0
		input  wire [7:0]  datab_1, // datab_1.datab_1
		input  wire [7:0]  datab_2, // datab_2.datab_2
		input  wire [7:0]  datab_3, // datab_3.datab_3
		output wire [25:0] result   //  result.result
	);

	mult_add_fix8bx16bx4_altera_mult_add_180_4l2tjzi mult_add_0 (
		.result  (result),  //  output,  width = 26,  result.result
		.dataa_0 (dataa_0), //   input,  width = 16, dataa_0.dataa_0
		.dataa_1 (dataa_1), //   input,  width = 16, dataa_1.dataa_1
		.dataa_2 (dataa_2), //   input,  width = 16, dataa_2.dataa_2
		.dataa_3 (dataa_3), //   input,  width = 16, dataa_3.dataa_3
		.datab_0 (datab_0), //   input,   width = 8, datab_0.datab_0
		.datab_1 (datab_1), //   input,   width = 8, datab_1.datab_1
		.datab_2 (datab_2), //   input,   width = 8, datab_2.datab_2
		.datab_3 (datab_3), //   input,   width = 8, datab_3.datab_3
		.clock0  (clock0)   //   input,   width = 1,  clock0.clock0
	);

endmodule
